-- ----------------------------------------------------
-- Engineer : <Sergio Mercado Nunez > ( <SM9276@RIT.EDU>)
--
-- Create Date : <10/20/24 >
-- Design Name : globals
-- Module Name : globals - package ( library )
-- Project Name : < GameBoy-VHDL >
--
-- Description :
-- ----------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
package globals is
    constant Z_flag : integer := 7;
    constant N_flag : integer := 6;
    constant H_flag : integer := 5;
    constant C_flag : integer := 4;
end;

